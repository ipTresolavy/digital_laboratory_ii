../../../exp1/simulation/controle_servo.vhd