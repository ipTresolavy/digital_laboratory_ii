../../../exp1/simulation/controle_servo_tb.vhd