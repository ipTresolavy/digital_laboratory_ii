../simulation/controle_servo_tb.vhd