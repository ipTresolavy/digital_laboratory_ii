../simulation/circuito_pwm_tb.vhd