../simulation/circuito_pwm.vhd