../simulation/controle_servo.vhd