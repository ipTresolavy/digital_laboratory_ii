../../../exp1/simulation/circuito_pwm_tb.vhd