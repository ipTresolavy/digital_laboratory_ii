../../../exp1/simulation/counter.vhd