../../../exp1/simulation/desafio.vhd