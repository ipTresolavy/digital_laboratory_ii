../../../exp1/simulation/circuito_pwm.vhd